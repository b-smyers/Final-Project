module LeftShifterTwoBits(ValueIn, ValueOut); // to calc. JumpAddr for J instruction
  input [25:0] ValueIn; // 26-bit input
  output [27:0] ValueOut; // 28-bit output

endmodule
