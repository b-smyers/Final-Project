module BEQAdder(ValueIn1, ValueIn2, ValueOut); // PC+4+Jumpaddr BEQ jump address
  input [31:0] ValueIn1, ValueIn2; // 32-bit inputs
  output [31:0] ValueOut; // sum of inputs

endmodule
