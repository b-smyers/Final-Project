module PCAdder(PCIn, PCOut);
  input [31:0] PCIn; // 32-bit address
  input [31:0] PCOut; // input incremented by 4

endmodule
